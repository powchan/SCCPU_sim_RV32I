library verilog;
use verilog.vl_types.all;
entity sccomp is
    port(
        clk             : in     vl_logic;
        rstn            : in     vl_logic
    );
end sccomp;
